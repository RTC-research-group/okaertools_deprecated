--
--	Package File Template
--
--	Purpose: This package defines supplemental types, subtypes, 
--		 constants, and functions 
--
--   To use any of the example code shown below, uncomment the lines and modify as necessary
--

library IEEE;
use IEEE.STD_LOGIC_1164.all;

package okt_imu_pkg is

end okt_imu_pkg;

package body okt_imu_pkg is
 
end okt_imu_pkg;
